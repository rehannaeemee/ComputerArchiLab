module testbench


initial begin

	test_PC;
	test_IM;
	test_ALU;
	test_RegFile;
	test_DM;
	test_IG;
	test_adders;

end

endmodule